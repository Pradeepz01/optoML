module pipeline_reg #(
    parameter DATA_WIDTH = 32
)(
    input  logic                   clk,
    input  logic                   rst_n,

    // Input interface
    input  logic                   in_valid,
    output logic                   in_ready,
    input  logic [DATA_WIDTH-1:0]  in_data,

    // Output interface
    output logic                   out_valid,
    input  logic                   out_ready,
    output logic [DATA_WIDTH-1:0]  out_data
);

    // Internal storage
    logic [DATA_WIDTH-1:0] data_reg;
    logic                  valid_reg;

    // Ready when storage is empty OR output is consuming data
    assign in_ready = ~valid_reg || (out_ready && out_valid);

    // Output assignments
    assign out_valid = valid_reg;
    assign out_data  = data_reg;

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            valid_reg <= 1'b0;
        end
        else begin
            // Accept new data
            if (in_valid && in_ready) begin
                data_reg  <= in_data;
                valid_reg <= 1'b1;
            end
            // Output consumed with no new input
            else if (out_ready && out_valid) begin
                valid_reg <= 1'b0;
            end
        end
    end

endmodule
